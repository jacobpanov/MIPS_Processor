// Jacob Panov
// This module implements a controller for a simple CPU architecture.
// controller.v

`include "definitions.v"

module controller ()