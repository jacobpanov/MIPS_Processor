// Jacob Panov
//
// top.sv

`include "definitions.sv"

